module (input logic A,B,C,D,E,F,
			output logic H,I,J,K,L,M,N);
			
		assign H = (A & B) | (A & C);
		
		
endmodule