-- Restador completo de 4 std_logics
library IEEE;
use IEEE.std_logic_1164.all;

 
entity rest4std_logic is
	port(A,B: in std_logic_vector(3 downto 0);-- 4 entradas 
			Bin : in std_logic;
			Sf: out std_logic_vector(4 downto 0));-- 5 salidas (1 borrow y 4 de resultado)
end entity;


architecture structural of rest4std_logic is
	Signal Borrow: std_logic_vector(2 downto 0);-- Borrows
	--Declaración de componentes
	component rest1std_logic is
		port(Ai,Bi,Bin: in std_logic;
				S,Bout: out std_logic);
	end component rest1std_logic;
	
	begin
	--Sf(0),..,sf(3) = resultado de la resta
	--sf(4) = Borrow de salida
		rest0: rest1std_logic
			port map(Ai=>A(0),Bi=>B(0),Bin=>Bin,S=>Sf(0),Bout=>Borrow(0));
		rest1: rest1std_logic
			port map(Ai=>A(1),Bi=>B(1),Bin=>Borrow(0),S=>Sf(1),Bout=>Borrow(1));
		rest2: rest1std_logic
			port map(Ai=>A(2),Bi=>B(2),Bin=>Borrow(1),S=>Sf(2),Bout=>Borrow(2));
		rest3: rest1std_logic
			port map(Ai=>A(3),Bi=>B(3),Bin=>Borrow(2),S=>Sf(3),Bout=>Sf(4));	
	
end architecture;